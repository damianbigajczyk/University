library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CNT10 is
    Port ( RESET : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           C : out  STD_LOGIC;
           Q : out  STD_LOGIC_VECTOR (3 downto 0));
end CNT10;

architecture Behavioral of CNT10 is

begin


end Behavioral;

