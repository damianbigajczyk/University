library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Detektor_sekwencji_1010 is
    Port ( I : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           RESET : in  STD_LOGIC;
           O : out  STD_LOGIC);
end Detektor_sekwencji_1010;

architecture Behavioral of Detektor_sekwencji_1010 is

begin


end Behavioral;

