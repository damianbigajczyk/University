`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:47:16 03/16/2019 
// Design Name: 
// Module Name:    BINTO7SEG 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BINTO7SEG(
    input [3:0] BIN,
    input DP,
    input EN,
    output [7:0] SEG
    );


endmodule
